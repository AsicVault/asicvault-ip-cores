reg [P_UC_WIDTH-1:0] testcode[] = '{
14'h0000, //    0: LDW 0
14'h0081, //    1: ADDW 1
14'h187F, //    2: STW 63
14'h00C0, //    3: ADDX2 0
14'h187E, //    4: STW 62
14'h0104, //    5: SUBW 4
14'h01C0, //    6: SHRW
14'h1855, //    7: STW 21
14'h013E, //    8: SUBW 62
14'h1854, //    9: STW 20
14'h0000, //   10: LDW 0
14'h0503, //   11: SUBW 3 KEEP_W
14'h240B, //   12: TSS CARRY
14'h3067, //   13: JUMP TEST1_ERROR1 = 116
14'h2402, //   14: TSC ZERO
14'h3066, //   15: JUMP TEST1_ERROR2 = 117
14'h0100, //   16: SUBW 0
14'h2403, //   17: TSS ZERO
14'h3064, //   18: JUMP TEST1_ERROR3 = 118
14'h240A, //   19: TSC CARRY
14'h3063, //   20: JUMP TEST1_ERROR4 = 119
14'h3002, //   21: JUMP +2
14'h2000, //   22: NOP
14'h1845, //   23: STW 5
14'h0001, //   24: LDW 1
14'h0200, //   25: MUL_PUSH 0
14'h1ABD, //   26: MUL_STH 61
14'h1E7C, //   27: MUL_POP 60 keep_w
14'h0202, //   28: MUL_PUSH 2
14'h0203, //   29: MUL_PUSH 3
14'h1A9F, //   30: MUL_STH 31
14'h1E5E, //   31: MUL_POP 30 keep_w
14'h1AA1, //   32: MUL_STH 33
14'h1E60, //   33: MUL_POP 32 keep_w
14'h3008, //   34: jump JTEST1 = 42
14'h0004, //   35: LDW 4
14'h0101, //   36: SUBW 1
14'h0101, //   37: SUBW 1
14'h184B, //   38: STW 11
14'h2407, //   39: STOP 
14'h0000, //   40: LDW 0
14'h0001, //   41: LDW 1
14'h0003, //   42: LDW 3
14'h0100, //   43: SUBW 0
14'h184A, //   44: STW 10
14'h3FF7, //   45: go JTEST2 = 36 
14'h0000, //   46: LDW 0
14'h0186, //   47: HFPRIM 6
14'h0186, //   48: HFPRIM 6
14'h1847, //   49: STW 7
14'h0001, //   50: LDW 1
14'h0186, //   51: HFPRIM 6
14'h0186, //   52: HFPRIM 6
14'h1848, //   53: STW 8
14'h0002, //   54: LDW 2
14'h0186, //   55: HFPRIM 6
14'h0186, //   56: HFPRIM 6
14'h1849, //   57: STW 9
14'h2407, //   58: STOP 
14'h000A, //   59: LDW 10
14'h020B, //   60: MUL_PUSH 11
14'h000C, //   61: LDW 12
14'h020D, //   62: MUL_PUSH 13
14'h1A8F, //   63: MUL_STH 15
14'h1A4E, //   64: MUL_POP 14
14'h1A91, //   65: MUL_STH 17
14'h1A50, //   66: MUL_POP 16
14'h2407, //   67: STOP 
14'h2809, //   68: LOOPINIT 9
14'h001E, //   69: LDW 30
14'h2433, //   70: TSS W0
14'h3003, //   71: jump +3
14'h001F, //   72: LDW 31
14'h02E0, //   73: MUL_PUSH_CPRIME 32
14'h001F, //   74: LDW 31
14'h02DF, //   75: MUL_PUSH_CPRIME 31
14'h2442, //   76: TSC LAST
14'h1B60, //   77: CPRIME_POP 32
14'h1B5F, //   78: CPRIME_POP 31
14'h001E, //   79: LDW 30
14'h01C0, //   80: SHRW
14'h185E, //   81: STW 30
14'h243B, //   82: TSS LOOPDONE
14'h3FF3, //   83: jump BINV_LOOP1 = 70 
14'h2815, //   84: LOOPINIT 21
14'h001F, //   85: LDW 31
14'h02DF, //   86: MUL_PUSH_CPRIME 31
14'h02E0, //   87: MUL_PUSH_CPRIME 32
14'h243A, //   88: TSC LOOPDONE
14'h3006, //   89: jump BINV_LOOP_OUT1 = 95
14'h1B5F, //   90: CPRIME_POP 31
14'h1F60, //   91: CPRIME_POP 32 keep_w
14'h02DF, //   92: MUL_PUSH_CPRIME 31
14'h02E0, //   93: MUL_PUSH_CPRIME 32
14'h3FFA, //   94: jump BINV_LOOP_P1 = 88 
14'h1B5F, //   95: CPRIME_POP 31
14'h1F60, //   96: CPRIME_POP 32 keep_w
14'h02DF, //   97: MUL_PUSH_CPRIME 31
14'h1B5F, //   98: CPRIME_POP 31
14'h28DE, //   99: LOOPINIT 222
14'h02DF, //  100: MUL_PUSH_CPRIME 31
14'h02E0, //  101: MUL_PUSH_CPRIME 32
14'h243A, //  102: TSC LOOPDONE
14'h3006, //  103: jump BINV_FINISH = 109
14'h1B5F, //  104: CPRIME_POP 31
14'h1F60, //  105: CPRIME_POP 32 keep_w
14'h02DF, //  106: MUL_PUSH_CPRIME 31
14'h02E0, //  107: MUL_PUSH_CPRIME 32
14'h3FFA, //  108: jump BINV_LOOP2 = 102 
14'h1B5F, //  109: CPRIME_POP 31
14'h1B60, //  110: CPRIME_POP 32
14'h2407, //  111: STOP 
14'h000C, //  112: LDW 12
14'h030D, //  113: CPRIME_PUSH 13
14'h1B4E, //  114: CPRIME_POP 14
14'h2407, //  115: STOP 
14'h2407, //  116: STOP 
14'h2407, //  117: STOP 
14'h2407, //  118: STOP 
14'h2407  //  119: STOP 
};
//PROC Start positions:
const reg [P_UC_WIDTH-1:0] PRIME_ONLY_TEST = 14'h0070;
const reg [P_UC_WIDTH-1:0] BINV_TEST = 14'h0044;
const reg [P_UC_WIDTH-1:0] TEST3 = 14'h003B;
const reg [P_UC_WIDTH-1:0] TEST2 = 14'h002E;
const reg [P_UC_WIDTH-1:0] TEST1 = 14'h0000;

